library verilog;
use verilog.vl_types.all;
entity cu_vlg_vec_tst is
end cu_vlg_vec_tst;
