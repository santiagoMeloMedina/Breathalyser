library verilog;
use verilog.vl_types.all;
entity pc_memory_control_tb_vlg_vec_tst is
end pc_memory_control_tb_vlg_vec_tst;
