library verilog;
use verilog.vl_types.all;
entity pc_memory_control_tb_vlg_sample_tst is
    port(
        reloj           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end pc_memory_control_tb_vlg_sample_tst;
