library verilog;
use verilog.vl_types.all;
entity arm_vlg_vec_tst is
end arm_vlg_vec_tst;
