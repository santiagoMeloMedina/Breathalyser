library verilog;
use verilog.vl_types.all;
entity am_vlg_vec_tst is
end am_vlg_vec_tst;
